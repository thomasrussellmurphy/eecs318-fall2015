// Thomas Russell Murphy (trm70)
// EECS 318 Fall 2015
// The implementation a full-adder with a 10 unit gate delay
// Will be used for implementing a ripple-carry adder

`timescale 1 ns / 1 ps

module adder(
         input A, B, Ci,
         output S, Co
       );

wire ABsum;
wire ABcarry, Ccarry;

// Compute the sum
xor #10 ( ABSum, A, B );
xor #10 ( S, Ci, ABsum );

// Compute the ripple-carry
and #10 ( Ccarry, ABsum, Ci );
and #10 ( ABcarry, A, B );
or #10 ( Co, Ccarry, ABcarry );

endmodule
