-- Thomas Russell Murphy (trm70)
-- EECS 318 Fall 2015
-- Generic width ripple-carry adder

library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.STD_LOGIC_ARITH.ALL;
  use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity csa_10_8 is
  port (
  a : in std_logic_vector(7 downto 0);
  b : in std_logic_vector(7 downto 0);
  c : in std_logic_vector(7 downto 0);
  d : in std_logic_vector(7 downto 0);
  e : in std_logic_vector(7 downto 0);
  f : in std_logic_vector(7 downto 0);
  g : in std_logic_vector(7 downto 0);
  h : in std_logic_vector(7 downto 0);
  i : in std_logic_vector(7 downto 0);
  j : in std_logic_vector(7 downto 0);
  z : out std_logic_vector(11 downto 0) );

end csa_10_8;

architecture RTL of adder_rc is
  -- Signals

  -- Components
begin
  -- Layer 1
  -- Layer 2
  -- Layer 3
  -- Layer 4
  -- Layer 5
  -- Final adder
end RTL;
